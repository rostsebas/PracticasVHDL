----------------------------------------------------------------------------------
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity Multiplexacion is
	port(
		clk : in	std_logic;
		canal1, canal2 : in std_logic
	);
end Multiplexacion;

architecture Behavioral of Multiplexacion is

begin


end Behavioral;

